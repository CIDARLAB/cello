module structuralAND(output out, input inA, inB);

   and (out, inA, inB);
   
endmodule

