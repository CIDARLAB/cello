
        2'b11: {out1} = 1'b1;
      endcase
    end
endmodule
