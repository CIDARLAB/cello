module structuralNOT(output out, input inA);

   not (out, inA);
   
endmodule

